// -----------------------------------------------------------------------------
// Copyright (c) 2020 All rights reserved
// -----------------------------------------------------------------------------
// Author   : Shubhasini D (shubhasinid@gmail.com)
// File     : 43_gnd.v
// Create   : 2020-08-30 15:52:15
// Revise   : 2020-08-30 15:52:16
// Comments :
// -----------------------------------------------------------------------------


module top_module (
	output out
);
	assign out = 1'b0;
endmodule
