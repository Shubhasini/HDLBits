// -----------------------------------------------------------------------------
// Copyright (c) 2020 All rights reserved
// -----------------------------------------------------------------------------
// Author   : Shubhasini D (shubhasinid@gmail.com)
// File     : 42_wire.v
// Create   : 2020-08-30 15:52:08
// Revise   : 2020-08-30 15:52:09
// Comments :
// -----------------------------------------------------------------------------

module top_module (
	input  in ,
	output out
);
	assign out = in;
endmodule
