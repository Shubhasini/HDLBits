// -----------------------------------------------------------------------------
// Copyright (c) 2020 All rights reserved
// -----------------------------------------------------------------------------
// Author   : Shubhasini D (shubhasinid@gmail.com)
// File     : 77_kmap7.v
// Create   : 2020-08-30 17:23:00
// Revise   : 2020-08-30 17:27:13
// Comments :
// -----------------------------------------------------------------------------

module top_module (
	input  [4:1] x,
	output       f
);
	assign f = (~x[2] & ~x[4]) | (~x[1] & x[3]) |(x[2] & x[3] & x[4]);
endmodule
