// -----------------------------------------------------------------------------
// Copyright (c) 2020 All rights reserved
// -----------------------------------------------------------------------------
// Author                 : Shubhasini D (shubhasinid@gmail.com)
// File                   : 153_review2015_fsmshift.v
// Create                 : 2020-11-18 20:16:38
// Revision               : 2020-11-18 20:16:39
// url of que.            : https://hdlbits.01xz.net/wiki/Exams/review2015_fsmshift
// Description            :
//
// -----------------------------------------------------------------------------

module top_module (
    input clk,
    input reset,      // Synchronous reset
    output shift_ena);

endmodule
