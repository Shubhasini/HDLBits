//simple_wire.v

module top_module (
	input  in ,
	output out
);
	assign out = in; //connecting through wire
endmodule
