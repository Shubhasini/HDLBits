//replication.v
module top_module (
	input  [ 7:0] in ,
	output [31:0] out
);
//
// Concatenate two things together:
// 1: {in[7]} repeated 24 times (24 bits)
// 2: in[7:0] (8 bits)
	assign out[31:0] = { {24{in[7]}},in[7:0] };

endmodule
