// -----------------------------------------------------------------------------
// Copyright (c) 2020 All rights reserved
// -----------------------------------------------------------------------------
// Author           : Shubhasini D (shubhasinid@gmail.com)
// File             : 112_2014_q4b.v
// Create           : 2020-09-08 20:13:05
// Revision         : 2020-09-08 20:13:16
// Description      :
// 
// -----------------------------------------------------------------------------

module top_module (
    input [3:0] SW,
    input [3:0] KEY,
    output [3:0] LEDR
); //

endmodule

module MUXDFF (...);

endmodule
