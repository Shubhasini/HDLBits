// -----------------------------------------------------------------------------
// Copyright (c) 2020 All rights reserved
// -----------------------------------------------------------------------------
// Author   : Shubhasini D (shubhasinid@gmail.com)
// File     : 1_wire.v
// Create   : 2020-08-30 15:45:20
// Revise   : 2020-08-30 15:45:21
// Comments :
// -----------------------------------------------------------------------------


module top_module (
	input  in ,
	output out
);
	assign out = in; //connecting through wire
endmodule
